// Generate a square wave on a pin (not LED)

module square_wave # (

) (
    input 
);

endmodule
