// The following registers are "buckets" that hold the current color state.
// At the beginning of each "shift" cycle (of which there are 6 * SHIFT_COLORS),
// this_shift_p/f registers are assigned values that sum to 32. The distribution
// of those values depends on how much of a certain color is desired. 
// "p" and "f" refer to past and future, so if RED is the past color and MAGENTA the future, 
// and we desire a color that is more red than magenta, then the value assigned to this_shift_p
// will be larger than this_shift_f. The "prev_" variables simply keep track of the previous shift color
// so we can perform a smooth transition across the rainbow.
// On each shift_clk, one of this_shift_p/f is decremented if it is not empty. 
// The result is a rapid toggle between two neighboring colors that the human eye
// averages to make a single color between the two. By increasing the amount of "future" color 
// on each shift cycle, we circularly transition between colors.

module rainbow_led (
    input clk,
    input button_a,
    input button_b,

    output reg [2:0] led
);

wire rst = !button_a;

// base colors
localparam WHITE    = 3'b000;
localparam MAGENTA  = 3'b001;
localparam YELLOW   = 3'b010;
localparam RED      = 3'b011;
localparam CYAN     = 3'b100;
localparam BLUE     = 3'b101;
localparam GREEN    = 3'b110;
localparam OFF      = 3'b111;

localparam N_BASE_COLORS        = 6;    // 6 because WHITE/OFF are non-colors, in this case
localparam N_M_COLORS_PER_BASE  = 3;    // num minor colors between eash base color
localparam N_MINOR_COLORS       = N_M_COLORS_PER_BASE * N_BASE_COLORS;  // total num minor colors

localparam TICKS_PER_SEC        = 24_000_000;                       // system clk speed
localparam RAINBOW_SECS         = 10;                               // seconds per rainbow cycle
localparam RAINBOW_TICKS        = TICKS_PER_SEC * RAINBOW_SECS;     // clk ticks per rainbow cycle

localparam MINOR_COLOR_TICKS = RAINBOW_TICKS / N_MINOR_COLORS;   // ticks per minor color
localparam BLUR_TICKS = MINOR_COLOR_TICKS / N_M_COLORS_PER_BASE; // number of clk ticks in each shift slot

// drive blur color shift
reg [$clog2(BLUR_TICKS)-1:0] blur_clk_cnt = 0;
wire shift_blur_color = (blur_clk_cnt == BLUR_TICKS);
always @(posedge clk) begin
    if (shift_blur_color) begin
        blur_clk_cnt <= 0;
    end else begin
        blur_clk_cnt <= blur_clk_cnt + 1;
    end
end

// drive minor color shift
reg [$clog2(MINOR_COLOR_TICKS)-1:0] minor_clk_cnt = 0;
wire shift_minor_color = (minor_clk_cnt == MINOR_COLOR_TICKS);
always @(posedge clk) begin
    if (shift_minor_color) begin
        minor_clk_cnt <= 0;
    end else begin
        minor_clk_cnt <= minor_clk_cnt + 1;
    end
end

// drive base color shift
reg [$clog2(N_M_COLORS_PER_BASE)-1:0] base_clk_cnt = 0;
wire shift_base_color = (base_clk_cnt == N_M_COLORS_PER_BASE);
always @(posedge shift_minor_color) begin
    if (shift_base_color) begin
        base_clk_cnt <= 0;
    end else begin
        base_clk_cnt <= base_clk_cnt + 1;
    end
end

// shift base color
always @(posedge shift_base_color) begin
    past_base_color     <= future_base_color;
    future_base_color   <= past_base_color;
end

// reset to next minor color or pick current blur color
reg [2:0] past_base_color    = RED;
reg [2:0] future_base_color  = ~RED;

localparam W = $clog2(N_M_COLORS_PER_BASE)-1;
reg [W:0] last_past_blur_col = 0;
reg [W:0] last_fut_blur_col  = 0;
reg [W:0] this_past_blur_col = N_M_COLORS_PER_BASE;
reg [W:0] this_fut_blur_col  = 0;

always @(shift_minor_color) begin
    this_past_blur_col  <= last_past_blur_col - 1;
    this_fut_blur_col   <= last_fut_blur_col + 1;
    
    last_past_blur_col  <= this_past_blur_col;
    last_fut_blur_col   <= this_fut_blur_col;
    
    this_past_blur_col  <= this_past_blur_col - 1;
    this_fut_blur_col   <= this_fut_blur_col - 1;
end

wire p_empty = (this_past_blur_col  == 0);
wire f_empty = (this_fut_blur_col   == 0);

always @(posedge shift_blur_color) begin
    if (!p_empty) begin
        led <= past_base_color;
    end else if (!f_empty) begin
        led <= future_base_color;
    end else begin
        led <= GREEN;
    end
end    
endmodule